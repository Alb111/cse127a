
package config_pkg;

  // define structs and enums needed for design
  parameter int ADDR_WIDTH = 32;
  parameter int MEM_WIDTH = 32;
  parameter int CountWidth = 8;

endpackage
