module mem_ctrl import config_pkg::*; #(
) (
    input  logic clk_i,
    input  logic rst_ni,
    output logic led_o
);

endmodule
